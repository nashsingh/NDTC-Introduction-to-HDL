LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Lab2_Part1 IS
PORT (SW0: 	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		SW1: 	IN STD_LOGIC_VECTOR(7 DOWNTO 4);
		HEX0: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX1: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX2: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX3: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
		
		END Lab2_Part1;
		
		ARCHITECTURE Behavior OF Lab2_Part1 IS 
		BEGIN 
		
		HEX0 <= "1000000" WHEN SW0 = "0000" ELSE
				  "1111001" WHEN SW0 = "0001" ELSE
				  "0100100" WHEN SW0 = "0010" ELSE
				  "0110000" WHEN SW0 = "0011" ELSE
				  "0011001" WHEN SW0 = "0100" ELSE
				  "0010010" WHEN SW0 = "0101" ELSE
				  "0000010" WHEN SW0 = "0110" ELSE
				  "1011000" WHEN SW0 = "0111" ELSE
				  "0000000" WHEN SW0 = "1000" ELSE
				  "0011000" WHEN SW0 = "1001" ELSE
				  "1111111" ;
				  
		HEX1 <= "1000000" WHEN SW1 = "0000" ELSE
				  "1111001" WHEN SW1 = "0001" ELSE
				  "0100100" WHEN SW1 = "0010" ELSE
				  "0110000" WHEN SW1 = "0011" ELSE
				  "0011001" WHEN SW1 = "0100" ELSE
				  "0010010" WHEN SW1 = "0101" ELSE
				  "0000010" WHEN SW1 = "0110" ELSE
				  "1011000" WHEN SW1 = "0111" ELSE
				  "0000000" WHEN SW1 = "1000" ELSE
				  "0011000" WHEN SW0 = "1001" ELSE
				  "1111111" ;
				  
		HEX2 <= "1111111";
		
		HEX3 <= "1111111";
				  
				  END Behavior;
				  
				 